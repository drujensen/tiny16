`timescale 1ns/1ns

module tiny16_tb;

endmodule
